library IEEE;
use IEEE.STD_LOGIC_1164.all;

-- notes Drawing 
entity NotesDrwaings is
port 	(
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoordY	: in integer;
		offset 		: in integer;
		mVGA_RGB    : out std_logic_vector(7 downto 0);
		soul_request	: out std_logic;
		drawing_requests	: out std_logic_vector(17 downto 0)
	);
end NotesDrwaings;

architecture behav of NotesDrwaings is 

--soul size
constant soul_X_size : integer := 45;
constant soul_Y_size : integer := 87;
--note size
constant note_X_size : integer := 25;
constant note_Y_size : integer := 60;

type object_form is array (0 to soul_Y_size - 1 , 0 to soul_X_size - 1) of std_logic;
--the soul image
constant soul : object_form := (
("000000000000000000000000111000000000000000000"),
("000000000000000000000001111100000000000000000"),
("000000000000000000000011111110000000000000000"),
("000000000000000000000111111110000000000000000"),
("000000000000000000000111111110000000000000000"),
("000000000000000000001111111111000000000000000"),
("000000000000000000001111111111000000000000000"),
("000000000000000000011111111111000000000000000"),
("000000000000000000011111100011000000000000000"),
("000000000000000000011111000011100000000000000"),
("000000000000000000011110000001100000000000000"),
("000000000000000000011110000001100000000000000"),
("000000000000000000111100000001100000000000000"),
("000000000000000000111100000001100000000000000"),
("000000000000000000111000000011100000000000000"),
("000000000000000000111000000011100000000000000"),
("000000000000000000111000000011100000000000000"),
("000000000000000000111000000111100000000000000"),
("000000000000000000011000000111100000000000000"),
("000000000000000000011000001111000000000000000"),
("000000000000000000011000011111000000000000000"),
("000000000000000000011000011111000000000000000"),
("000000000000000000011000111111000000000000000"),
("000000000000000000011001111110000000000000000"),
("000000000000000000001011111110000000000000000"),
("000000000000000000001111111110000000000000000"),
("000000000000000000001111111100000000000000000"),
("000000000000000000011111111100000000000000000"),
("000000000000000000111111111000000000000000000"),
("000000000000000001111111110000000000000000000"),
("000000000000000011111111110000000000000000000"),
("000000000000000111111111100000000000000000000"),
("000000000000000111111111000000000000000000000"),
("000000000000001111111110000000000000000000000"),
("000000000000011111111110000000000000000000000"),
("000000000000111111111110000000000000000000000"),
("000000000001111111110010000000000000000000000"),
("000000000011111111100011000000000000000000000"),
("000000000011111111000011000000000000000000000"),
("000000000111111110000011000000000000000000000"),
("000000000111111000000001000000000000000000000"),
("000000001111111000000001000000000000000000000"),
("000000001111110000000001111111000000000000000"),
("000000011111100000000111111111110000000000000"),
("000000011111000000001111111111111000000000000"),
("000000011111000000011111111111111100000000000"),
("000000011110000000111111111111111110000000000"),
("000000011110000001111111111111111111000000000"),
("000000111110000001111110110001111111000000000"),
("000000111110000011111100110000111111100000000"),
("000000011100000011111000010000011111100000000"),
("000000011100000011110000011000001111100000000"),
("000000011100000011110000011000001111100000000"),
("000000011100000011110000011000000111100000000"),
("000000011110000011110000011000000111100000000"),
("000000001110000011110000001000000111100000000"),
("000000001110000001110000001100000111100000000"),
("000000001110000000110000001100000111100000000"),
("000000000111000000011000001100000111100000000"),
("000000000011000000001100001100000111000000000"),
("000000000011100000000110001100001111000000000"),
("000000000001110000000000000110011110000000000"),
("000000000000111000000000000110111100000000000"),
("000000000000011110000000000111111000000000000"),
("000000000000000111110000000111110000000000000"),
("000000000000000011111111111111000000000000000"),
("000000000000000000001111110111000000000000000"),
("000000000000000000000000000011000000000000000"),
("000000000000000000000000000011000000000000000"),
("000000000000000000000000000011000000000000000"),
("000000000000000000000000000011000000000000000"),
("000000000000000000000000000011000000000000000"),
("000000000000000000000000000001100000000000000"),
("000000000000000000100000000001100000000000000"),
("000000000000000011111100000001100000000000000"),
("000000000000000111111100000001100000000000000"),
("000000000000001111111110000001100000000000000"),
("000000000000001111111110000001100000000000000"),
("000000000000011111111110000001100000000000000"),
("000000000000011111111110000001100000000000000"),
("000000000000011111111100000001100000000000000"),
("000000000000011111111000000001100000000000000"),
("000000000000001111100000000011000000000000000"),
("000000000000000111100000000111000000000000000"),
("000000000000000011110000011110000000000000000"),
("000000000000000001111111111100000000000000000"),
("000000000000000000001111110000000000000000000")
);

type note_ram_array is array(0 to note_Y_size - 1 , 0 to note_X_size - 1) of std_logic;
-- array for the notes image
constant note1: note_ram_array :=(
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000111111100000"),
("0000000000001111111100000"),
("0000000000011111111100000"),
("0000000000111111111100000"),
("0000000000111111111100000"),
("0000000001111111111100000"),
("0000000001111111111100000"),
("0000000001111111111100000"),
("0000000011111111111100000"),
("0000000011111111111000000"),
("0000000011111111111000000"),
("0000000001111111110000000"),
("0000000001111111100000000"),
("0000000000111111000000000"),
("0000000000011100000000000"),
("0000000000000000000000000")
); 
constant note2: note_ram_array :=(
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000011111111100000"),
("0000000000111111111100000"),
("0000000011111110001100000"),
("0000000111111000001100000"),
("0000000111110000001100000"),
("0000001111100000001100000"),
("0000001111000000011100000"),
("0000011110000000111100000"),
("0000011100000000111100000"),
("0000011100000001111000000"),
("0000011000000011111000000"),
("0000001000001111110000000"),
("0000001000111111100000000"),
("0000001111111111000000000"),
("0000000111111100000000000"),
("0000000011111000000000000"),
("0000000000000000000000000")
);
constant note3: note_ram_array :=(
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000000000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000000000100000"),
("0000000000000001000100000"),
("0000000000001001000100000"),
("0000000000001001000100000"),
("0000000000001001100100000"),
("0000000000001111100100000"),
("0000000000011111000100000"),
("0000000000011001000100000"),
("0000000000001001000100000"),
("0000000000001001000100000"),
("0000000000001001100100000"),
("0000000000001111100100000"),
("0000000000011111100100000"),
("0000000000011101000100000"),
("0000000000001001000100000"),
("0000000000001001000100000"),
("0000000000001000000100000"),
("0000000000000000000100000"),
("0000000000000111111100000"),
("0000000000001111111100000"),
("0000000000011111111100000"),
("0000000000111111111100000"),
("0000000000111111111100000"),
("0000000001111111111100000"),
("0000000001111111111100000"),
("0000000001111111111100000"),
("0000000011111111111100000"),
("0000000011111111111000000"),
("0000000011111111111000000"),
("0000000001111111110000000"),
("0000000001111111100000000"),
("0000000000111111000000000"),
("0000000000011100000000000"),
("0000000000000000000000000")
);
--soul boundaries
signal bCoord_X : integer := 0;
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

--notes boundaries
signal note_X_Coord : integer := 0;
signal note_Y_Coord : integer := 0;
signal note_Y_Coord_Down : integer :=0 ;

signal note_drawing_X : std_logic := '0';
signal note_drawing_Y : std_logic := '0';
signal note_drawing_Y_Down : std_logic :='0' ;
--		
signal objectWestXboundary : integer;
constant SoulStartX : integer := 10;
constant SoulStartY : integer := 45;

signal oCoord_Y :integer;
signal oCoord_Y_Down : integer ;

begin

--fixed coord_Y after offset
oCoord_Y	<= oCoordY+offset-7 when (offset < 100) and (oCoord_X  >= 55) else oCoordY-7;

-- Calculate Soul boundaries
objectWestXboundary	<= soul_X_size+SoulStartX;


--calculating  x & y coordination for drawing the pictures
-- Signals drawing_X[Y] are active when objects coordinates are being crossed

--for soul
	drawing_X	<= '1' when  (oCoord_X  >= SoulStartX) and  (oCoord_X < objectWestXboundary) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= SoulStartY) and  (oCoord_Y  < 400) and ((oCoord_Y-SoulStartY)mod(120) < soul_Y_size) else '0';

	bCoord_X 	<= (oCoord_X - SoulStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (((oCoord_Y-SoulStartY)mod(120))mod(87)) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
--for notes
	note_drawing_X	<= '1' when  (oCoord_X  >= 55) and  (oCoord_X < 605) else '0';
    note_drawing_Y	<= '1' when  (oCoord_Y  >= 75) and (oCoord_Y  < 400) and ((oCoord_Y-75)mod(120) < note_Y_size) else '0';

	note_X_Coord 	<= ((oCoord_X-55)mod(25)) when ( note_drawing_X = '1' and  note_drawing_Y = '1'  ) else 0 ; 
	note_Y_Coord 	<= (((oCoord_Y-75)mod(120))mod(60)) when ( note_drawing_X = '1' and  note_drawing_Y = '1'  ) else 0 ; 

process ( RESETn, CLK) 		
   begin
   	mVGA_RGB <= x"00" ;	
	if RESETn = '0' then	
		drawing_requests <= (others => '0');
		soul_request <= '0';
		elsif CLK'event and CLK='1' then
			if offset = 100 then
				drawing_requests <= (others=>'0');
			else
				-- create the different pictures
				drawing_requests(0) <= note_drawing_X and note_drawing_Y and note1(note_Y_Coord , note_X_Coord) ;--C4 /A
				drawing_requests(1) <= note_drawing_X and note_drawing_Y and note2(note_Y_Coord , note_X_Coord) ;--
				drawing_requests(2) <= note_drawing_X and note_drawing_Y and note2(note_Y_Coord , note_X_Coord) ;
				drawing_requests(3) <= note_drawing_X and note_drawing_Y and note3(note_Y_Coord , note_X_Coord) ;
				drawing_requests(4) <= note_drawing_X and note_drawing_Y and note2(note_Y_Coord , note_X_Coord) ;
				drawing_requests(5) <= note_drawing_X and note_drawing_Y and note2(note_Y_Coord , note_X_Coord) ;
				drawing_requests(6) <= note_drawing_X and note_drawing_Y and note1(note_Y_Coord , note_X_Coord) ;
				drawing_requests(7) <= note_drawing_X and note_drawing_Y and note2(note_Y_Coord , note_X_Coord) ;
				drawing_requests(8) <= note_drawing_X and note_drawing_Y and note2(note_Y_Coord , note_X_Coord) ;
				drawing_requests(9) <= note_drawing_X and note_drawing_Y and note3(note_Y_Coord , note_X_Coord) ;
				drawing_requests(10) <= note_drawing_X and note_drawing_Y and note2(note_Y_Coord , note_X_Coord) ;	
				drawing_requests(11) <= note_drawing_X and note_drawing_Y and note2(note_Y_Coord , note_X_Coord) ;
				drawing_requests(12) <= note_drawing_X and note_drawing_Y and note1(note_Y_size - note_Y_Coord ,note_X_size - note_X_Coord) ;	
				drawing_requests(13) <= note_drawing_X and note_drawing_Y and note2(note_Y_size - note_Y_Coord ,note_X_size - note_X_Coord) ;
				drawing_requests(14) <= note_drawing_X and note_drawing_Y and note3(note_Y_size - note_Y_Coord ,note_X_size - note_X_Coord) ;		
				drawing_requests(15) <= note_drawing_X and note_drawing_Y and note2(note_Y_size - note_Y_Coord ,note_X_size - note_X_Coord) ;
				drawing_requests(16) <= note_drawing_X and note_drawing_Y and note2(note_Y_size - note_Y_Coord ,note_X_size - note_X_Coord) ;	
				drawing_requests(17) <= note_drawing_X and note_drawing_Y and note2(note_Y_size - note_Y_Coord ,note_X_size - note_X_Coord) ;
				
--- using the 3 basic  pictures we can create 17 differnet notes shapes 

				--add "-" to the do image		
				if note_Y_Coord=48 and (note_X_Coord>4 and note_X_Coord<22) then
					if note_X_Coord>5 then
						drawing_requests(0) <= '1';
						drawing_requests(1) <= '1';
						drawing_requests(2) <= '1';
					drawing_requests(3) <= '1';
					end if;
					drawing_requests(4) <= '1';
					drawing_requests(5) <= '1';

				end if;
				--draw full circle(4/4) by keeping only the circle from the image 
				if (note_Y_Coord<44  and note_Y_Coord>=0 )or (note_Y_Coord=44  and note_X_Coord=19) then
					drawing_requests(2) <= '0';
					drawing_requests(5) <= '0';
					drawing_requests(8) <= '0';
					drawing_requests(11) <= '0';
				end if;
				if (note_Y_size - note_Y_Coord<43  and note_Y_size - note_Y_Coord>=0 )or (note_Y_size - note_Y_Coord=44  and note_X_Coord=19) then
					drawing_requests(16) <= '0';
					drawing_requests(17) <= '0';
				end if;
									
				-- add the "#" to the image
				if note_Y_Coord<43  and note_Y_Coord>26 and note_X_Coord < 17 then
					drawing_requests(4) <= note_drawing_X and note_drawing_Y and note3(note_Y_Coord , note_X_Coord) ;	
					drawing_requests(5) <= note_drawing_X and note_drawing_Y and note3(note_Y_Coord , note_X_Coord) ;	
					drawing_requests(10) <= note_drawing_X and note_drawing_Y and note3(note_Y_Coord , note_X_Coord) ;	
					drawing_requests(11) <= note_drawing_X and note_drawing_Y and note3(note_Y_Coord , note_X_Coord) ;	
				end if;
				if note_Y_size - note_Y_Coord<45  and note_Y_size - note_Y_Coord>27 and note_X_Coord < 15 then
					drawing_requests(15) <= note_drawing_X and note_drawing_Y and note3(note_Y_size - note_Y_Coord ,note_X_size - note_X_Coord) ;
					if  note_X_Coord > 9 then
						drawing_requests(17) <= note_drawing_X and note_drawing_Y and note3(note_Y_size - note_Y_Coord ,note_X_size - note_X_Coord) ;
					end if;
				end if;
			end if;
			-- draw the soul image 
			soul_request <= drawing_X and drawing_Y and soul(bCoord_Y , bCoord_X)  ;
			
	end if;
  end process;
end behav;		
		
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 -- flute table --
entity FluteSound is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(7 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end FluteSound;

architecture arch of FluteSound is

type table_type is array(0 to 255) of std_logic_vector(7 downto 0);
signal flute_table : table_type;

begin

  SinTableTC_proc: process(RESET_N, CLK,ADDR)
    constant flute_table : table_type := (
X"00",
X"02",
X"05",
X"07",
X"0A",
X"0C",
X"0F",
X"11",
X"14",
X"16",
X"19",
X"1B",
X"1E",
X"21",
X"23",
X"26",
X"28",
X"2B",
X"2D",
X"30",
X"32",
X"35",
X"37",
X"3A",
X"3C",
X"3F",
X"42",
X"44",
X"47",
X"49",
X"4C",
X"4E",
X"51",
X"53",
X"56",
X"58",
X"5B",
X"5D",
X"60",
X"63",
X"65",
X"68",
X"6A",
X"6D",
X"6F",
X"72",
X"74",
X"77",
X"79",
X"7C",
X"7F",
X"7F",
X"7D",
X"7C",
X"7B",
X"7A",
X"79",
X"78",
X"77",
X"76",
X"75",
X"74",
X"73",
X"72",
X"71",
X"70",
X"6F",
X"6E",
X"6D",
X"6C",
X"6B",
X"6A",
X"69",
X"68",
X"67",
X"66",
X"65",
X"64",
X"63",
X"62",
X"61",
X"60",
X"5F",
X"5E",
X"5D",
X"5B",
X"5A",
X"59",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"58",
X"57",
X"56",
X"55",
X"54",
X"53",
X"52",
X"51",
X"51",
X"50",
X"4F",
X"4E",
X"4D",
X"4C",
X"4B",
X"4A",
X"4A",
X"49",
X"48",
X"47",
X"46",
X"45",
X"44",
X"43",
X"43",
X"42",
X"41",
X"40",
X"3F",
X"3E",
X"3D",
X"3D",
X"3C",
X"3B",
X"3A",
X"39",
X"38",
X"37",
X"36",
X"36",
X"35",
X"34",
X"33",
X"32",
X"31",
X"30",
X"2F",
X"2F",
X"2E",
X"2D",
X"2C",
X"2B",
X"2A",
X"29",
X"28",
X"28",
X"27",
X"26",
X"25",
X"24",
X"23",
X"22",
X"21",
X"21",
X"20",
X"1F",
X"1E",
X"1D",
X"1C",
X"1B",
X"1B",
X"1A",
X"19",
X"18",
X"17",
X"16",
X"15",
X"14",
X"14",
X"13",
X"12",
X"11",
X"10",
X"0F",
X"0E",
X"0D",
X"0D",
X"0C",
X"0B",
X"0A",
X"09",
X"08",
X"07",
X"06",
X"06",
X"05",
X"04",
X"03",
X"02",
X"01",
X"00",
X"00"
  );

  begin

    if (RESET_N='0') then
      Q <= flute_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= flute_table(to_integer(unsigned(ADDR)));
      else
		Q <= flute_table(0);
	end if;
    end if;
  end process;
end arch;
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;

--drawing the background 

entity back_ground_draw is
	port(
		CLK  : in std_logic;
		RESETn	: in std_logic;
		oCoord_X 		: in integer;
		oCoord_Y 		: in integer;
		recording		: in std_logic;
		play			: in std_logic;
		mVGA_RGB	      : out std_logic_vector(7 downto 0) --	,  //	VGA Red[9:0]
	);
end back_ground_draw;

architecture behav of back_ground_draw is 

signal mVGA_R	: std_logic_vector(2 downto 0); --	,	 			//	VGA Red[9:0]
signal mVGA_G	: std_logic_vector(2 downto 0); --	,	 			//	VGA Green[9:0]
signal mVGA_B	:  std_logic_vector(1 downto 0); --	,  				//	VGA Blue[9:0]

---- drawing the lines----

--lines start
constant start : integer := 60;
--offset between each line
constant offset : integer := 15;
--distance between every 5 lines
constant dist : integer := 60;
 
 
---- drawing the welcome image ----

--size
constant welcome_X_size : integer := 283;
constant welcome_Y_size : integer :=27;

--object start
signal X_begin : integer := 180;
signal Y_begin : integer := 15 ;

signal bCoord_X : integer := 0;
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';


type Welcome_object is array (0 to welcome_Y_size - 1 , 0 to welcome_X_size - 1) of std_logic;
 constant welcome : Welcome_object := (
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011111111111"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000001110001110001111000000011100011111111111"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111100000001111000000000011111110001111000000001110001110001111000110011100011111111111"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000010000000001111110000000000000000111100100111100100001111000000001111111110001111000000001110001110001111100010011100011111111000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111000011100000000111100011111000111001000111111110000000000000001111100001111100110011111100100011111111110001111000000001110001110011111110010011100011100000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111001001111000011100000000111100111111000111000011111111110000000000000001111100001111100110011111100100111110000000001110011011001110001110011111110000011100011100000000"),
("0000000000000000000000000000000000000000000011110001110010000111111100110011110001001111000000000000000000000001111000001111100011100000000111101111110000111000011111100000000000000000001111110011111100100111111100000111100000000001110000000001110011110011111111000011100011100000000"),
("0000001100100011100000001111100000000011111111110001110000001111111100100011111001001111000000000000000000000011111100011111100011100000000111001111000000111000111100000000000000000000001111110011111100100111111110001111000000001001110000000011110011110011111111100011100011111111110"),
("0000111100100111110011001111100100000111111111110001110000111111111100100111111001001110000000000000000000000011111100011111100011100000000111001111001100111001111000000000000000000000011111111111111110001111011110001110000000000001111111111111110011110011110111110011100011111111110"),
("0000111110000111110010001111100110001111111111110001110001111110000000100111111001001110000000000000000000000011111110111111100011100000000111000111001100111001110000000000000000000000011111111111111110001111001110001110010000000001111111111111110011110011100111110011100011111111110"),
("0000111110001111110010011111110010011111000000000001110001111000000000001111111100001110000000000000000000000011111111111111100111100000000111000111100100111001110000000000000000000000011100111111011110001110001111011110000000000001111111111111110011110011100011111111100111100000000"),
("0001111110001111110010011111110000111100000000000001110011110000000011001111111100001110000000000000000000000011111111111111100111100000000111000111100100111011110000000000000000000000011100111110011110011110001111011110000000000001111000000011110011100011100001111111100111100000000"),
("0001111111011111110000111111110000111000000000000001110011100000000000011110011100001110000000000000000000000111101111110011100111100000000111000011110001111011110000000000000000000000111100111110001110011100001111001110000000001001110000000011110011100011100001111111100111100000000"),
("0001111111111111110000111101111001111001001111110001110111100000000000011110011110001110000000000000000000000111001111110011100111100000100111000011110001111011110000000000000000000000111100011100001110111111111111001111000000000001110011110011100011100011100100111111100111100000000"),
("0001111111111101110000111001111001110011001111110001110111100000000000011100011110001110000000000000000000000111000111100011110111100110000111001001111001111001110000000000000000000000111000011100001111111111111111101111100000000001110000000011100011100011100100011111100111111111111"),
("0011110111111101111001111001111001111011001111110011110111100000000000111100011110001110000000000000000000000111000111100011110111100010001111001001111001111001111000000000000000000000111001011001001111111111111111100111111111110011110000000011100011100011100110011111100111111111111"),
("0011110011111001111001110000111101111011001111110011110111100100000000111100001111001110010000000000000000001111000011000011110111110000011110000001111001111001111110000000000000000001111001001001001111111000000111100111111111110011110000000011100011100011100000001111100111111111111"),
("0011110011111001111011110000111101111001000011110011110011110000000001111111111111011110000000000000000000001111010011000011110011111101111110000011111001111000111111111110000000000001111001000001001111110000000011110001111111110011110000000011100011100011100000000111000000000000000"),
("0011100011110001111011111111111101111100000011110011110011111000000001111111111111011110000000000000000000001110010010011011110011111111111100001111111001111000011111111110000000000001111000000000001111110000010011110000011111100011100000000000000000000000000000000000000000000000000"),
("0111100001110001111111111111111110111110000011110011110011111110111011111111111111111111111111110000000000001110011000011011110001111111111000001111110001110010001111111110000000000001110000000000001111000000000011110010000000000000000000000000000000000000000000000000000000000000000"),
("0111100001100101111111111111111110111111111111110011110001111111111111110000000111111111111111110000000000011110000000000001110000011111100001001111100001110000000000000000000000000000000000000000001111000000000001111001000000000000000000000000000000000000000000000000000000000000000"),
("0111101100001101111111100000011110011111111111110011110100111111111111100000000111111111111111110000000000011110000000000001110010000000000000001110000000000000000000000000000000000000000000000000001111000000000001111000000000000000000000000000000000000000000000000000000000000000000"),
("0111001100001100111111000000001110000111111111110011110100001111111100100000000011111100000000000000000000000000000000000001111011000000000000000000000000000000000000000000000000000000000000000000000111000000000001110000000000000000000000000000000000000000000000000000000000000000000"),
("1111000000000100111110000001001111000001111111100000000000000000000000000000000011110000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("1111000000000000111100000000001111000000000011100000000000000000000000000000000011110010000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000111100000000001111001100000011100100000000000000000000000000000011110000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000111100000000000111100000000011100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);

---- drawing record image----

--record size
constant record_X_size : integer := 15;
constant record_Y_size : integer :=15;

--object start
signal X2_begin : integer := 150;
signal Y2_begin : integer := 400 ;

signal bCoord_X2 : integer := 0;
signal bCoord_Y2 : integer := 0;

signal drawing_X2 : std_logic := '0';
signal drawing_Y2 : std_logic := '0';


type record_object is array (0 to record_Y_size - 1 , 0 to record_X_size - 1) of std_logic;
 constant recording_img : record_object := (
("000000000000000"),
("000011111110000"),
("000111111111000"),
("001111111111100"),
("011111111111110"),
("011111111111110"),
("011111111111110"),
("111111111111111"),
("011111111111110"),
("011111111111110"),
("011111111111110"),
("001111111111100"),
("000111111111000"),
("000011111110000"),
("000000000000000")
);

----- play image -----
--size
constant play_X_size : integer := 15;
constant play_Y_size : integer :=16;

--object start
signal X3_begin : integer := 150;
signal Y3_begin : integer := 430;

signal bCoord_X3 : integer := 0;
signal bCoord_Y3 : integer := 0;

signal drawing_X3 : std_logic := '0';
signal drawing_Y3: std_logic := '0';


type play_object is array (0 to play_Y_size - 1 , 0 to play_X_size - 1) of std_logic;
 constant play_img : play_object := (
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111"),
("111110000011111")
);

begin

--calculating  x & y coordination for drawing the pictures

	drawing_X	<= '1' when  (oCoord_X  >=X_begin) and  (oCoord_X < X_begin+welcome_X_size) else '0';
	drawing_Y	<= '1' when  (oCoord_Y  >= Y_begin)  and (oCoord_Y  < Y_begin+welcome_Y_size) else '0';
            
	bCoord_X   <=  (oCoord_X-X_begin) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y   <= (oCoord_Y-Y_begin) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
------
	drawing_X2	<= '1' when  (oCoord_X  >=X2_begin) and  (oCoord_X < X2_begin+record_X_size) else '0';
	drawing_Y2	<= '1' when  (oCoord_Y  >= Y2_begin)  and (oCoord_Y  < Y2_begin+record_Y_size) else '0';
            
	bCoord_X2   <=  (oCoord_X-X2_begin) when ( drawing_X2 = '1' and  drawing_Y2 = '1'  ) else 0 ; 
	bCoord_Y2   <= (oCoord_Y-Y2_begin) when ( drawing_X2 = '1' and  drawing_Y2 = '1'  ) else 0 ; 
	
-----

	drawing_X3	<= '1' when  (oCoord_X  >=X3_begin) and  (oCoord_X < X3_begin+play_X_size) else '0';
	drawing_Y3	<= '1' when  (oCoord_Y  >= Y3_begin)  and (oCoord_Y  < Y3_begin+play_X_size) else '0';
            
	bCoord_X3   <=  (oCoord_X - X3_begin) when ( drawing_X3 = '1' and  drawing_Y3 = '1'  ) else 0 ; 
	bCoord_Y3   <= (oCoord_Y - Y3_begin) when ( drawing_X3 = '1' and  drawing_Y3 = '1'  ) else 0 ; 

--- drawing the lines in the background
mVGA_R <= "000" when 
	(  oCoord_y = start or oCoord_y = start+offset or oCoord_y = start+2*offset or oCoord_y = start+3*offset or oCoord_y = start+4*offset
	or oCoord_y = start+2*dist or oCoord_y = start+offset+2*dist or oCoord_y = start+2*offset+2*dist or oCoord_y = start+3*offset+2*dist or oCoord_y = start+4*offset+2*dist
	or oCoord_y = start+4*dist or oCoord_y = start+offset+4*dist or oCoord_y = start+2*offset+4*dist or oCoord_y = start+3*offset+4*dist or oCoord_y = start+4*offset+4*dist)
	else "111" ;	
mVGA_G <= "000" when
	(  oCoord_y = start or oCoord_y = start+offset or oCoord_y = start+2*offset or oCoord_y = start+3*offset or oCoord_y = start+4*offset
	or oCoord_y = start+2*dist or oCoord_y = start+offset+2*dist or oCoord_y = start+2*offset+2*dist or oCoord_y = start+3*offset+2*dist or oCoord_y = start+4*offset+2*dist
	or oCoord_y = start+4*dist or oCoord_y = start+offset+4*dist or oCoord_y = start+2*offset+4*dist or oCoord_y = start+3*offset+4*dist or oCoord_y = start+4*offset+4*dist)
	else "111" ;	
mVGA_B <= "00" when
	(  oCoord_y = start or oCoord_y = start+offset or oCoord_y = start+2*offset or oCoord_y = start+3*offset or oCoord_y = start+4*offset
	or oCoord_y = start+2*dist or oCoord_y = start+offset+2*dist or oCoord_y = start+2*offset+2*dist or oCoord_y = start+3*offset+2*dist or oCoord_y = start+4*offset+2*dist
	or oCoord_y = start+4*dist or oCoord_y = start+offset+4*dist or oCoord_y = start+2*offset+4*dist or oCoord_y = start+3*offset+4*dist or oCoord_y = start+4*offset+4*dist)
	else "11";
process (RESETn, CLK) 
begin
	 	if RESETn = '0' then
			mVGA_RGB <= (others =>'0');
		elsif rising_edge(CLK) then
			if  drawing_X='1' and drawing_Y='1' and (welcome(bCoord_Y , bCoord_X) ='1')then 
				mVGA_RGB <=  x"6F" ;-- draw the headline title  
			elsif drawing_X2='1' and drawing_Y2='1' and (recording_img(bCoord_Y2 , bCoord_X2) ='1') and recording ='1' then
				mVGA_RGB <=  x"e1" ;-- if the game in record state , show the record icon 
			elsif drawing_X3='1' and drawing_Y3='1' and (play_img(bCoord_Y3 , bCoord_X3)) ='1' and play ='1' then
				mVGA_RGB <=  x"00";-- if the game in play state , show the play icon 
			else
				mVGA_RGB <= mVGA_R & mVGA_G &  mVGA_B ; -- regrouping the colors in one vector 
			end if;
		end if;
	end process;
end behav;		
library IEEE;
use IEEE.STD_LOGIC_1164.all;

--- drawing the instruments screen 
entity Pick_inst_Screen is
port 	(
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		flute_effect		: in std_logic;
		piano_effect		:in std_logic ;
		drop_effect 		: in std_logic;
		pitch_effect		: in std_logic;
		Notes_screen_request : in std_logic;
		mVGA_RGB    : out std_logic_vector(7 downto 0);
		Pick_inst_request	: out std_logic
	);
end Pick_inst_Screen;

architecture behav of Pick_inst_Screen is 
--flute size
constant flute_X_size : integer :=66;
constant flute_Y_size : integer :=18;

--object start
signal X_begin : integer := 20;
signal Y_begin : integer := 400;

signal bCoord_X : integer := 0;
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';


type flute_object is array (0 to flute_Y_size - 1 , 0 to flute_X_size - 1) of std_logic;
 constant flute: flute_object := (
("000000000000000000000000000000000000000000000000000000000111111111"),
("000000000000000000000000000000000000000001101111111111100111111111"),
("000000000000000000000000000000001100000001101111111111100111000000"),
("011000000000001111100111000000001100000001101100111000000110000000"),
("111000000011111111100111000000001100000001100000111000000110000000"),
("111000000011111111100111000000001100000001100000111000000111111100"),
("111000000011000000000110000000001100000001100000111000001111111100"),
("111000000011000000000110000000001100000011100000111000001111100000"),
("111000000011000000000110000000001100000011100000111000001110000000"),
("111000000011111110000110000000001100000011100000110000001110000000"),
("111000000111111110000110000000011100000011100000110000001111111111"),
("111000000111100000000110000000001110000111000000110000001111111111"),
("111000000111000000000110000000001111111110000000110000001111111111"),
("111000000111000000001111111111000111111100000000110000000000000000"),
("111001100111000000001111111111000011111000000000000000000000000000"),
("111001100111000000001111111111000000000000000000000000000000000000"),
("111011100111000000000000000000000000000000000000000000000000000000"),
("111000000000000000000000000000000000000000000000000000000000000000")
);



 ----- piano image
constant piano_X_size : integer :=68;
constant piano_Y_size : integer :=19;
--object start
signal X2_begin : integer := 150;
signal Y2_begin : integer := 400;
 
signal bCoord_X2 : integer := 0;
signal bCoord_Y2 : integer := 0;

signal drawing_X2 : std_logic := '0';
signal drawing_Y2 : std_logic := '0';

type piano_object is array (0 to piano_Y_size - 1 , 0 to piano_X_size - 1) of std_logic;
 constant piano : piano_object := (
("00000000000000000000000000000000000000000000000000000000000001111000"),
("00000000000000000000000000000000000000000000001000000110000111111110"),
("00000000000000000000000000000000100001110000111100000110001111111111"),
("00001111100000000001111111100001100001110000111100000110011100000111"),
("00111111111000000011111111110011100011111000111110000110011000000011"),
("01111111111100000011111001111011100011111000111111000110111000000011"),
("11110000011100000011100000111011100111011000111111100110110000000011"),
("00100000011100000011000000011011100110011100110011101110110000000011"),
("00000000001110000011000000111011001110011100110011111110111000000111"),
("00000000001100000011000001110011001110001100110001111110111100001110"),
("00000000011100000011111111100011001111111110110000111110011111111100"),
("00000000011100000011111111000011111111111110110000111110001111111000"),
("00000000111100000011100000000011111100001111110000011110000011100000"),
("00000011111000110011000000000011111000000111110000000000000000000000"),
("00000111110001110011000000000011000000000111000000000000000000000000"),
("00001111100001110011000000000000000000000111000000000000000000000000"),
("00111110000000000000000000000000000000000011000000000000000000000000"),
("01111111111100000000000000000000000000000000000000000000000000000000"),
("11111111111100000000000000000000000000000000000000000000000000000000")
);
----- drop image
constant drop_X_size : integer :=68;
constant drop_Y_size : integer :=19;

--object start
signal X3_begin : integer := 320;
signal Y3_begin : integer := 400;

signal bCoord_X3 : integer := 0;
signal bCoord_Y3 : integer := 0;

signal drawing_X3 : std_logic := '0';
signal drawing_Y3 : std_logic := '0';

type drop_object is array (0 to drop_Y_size - 1 , 0 to drop_X_size - 1) of std_logic;
 constant drop : drop_object := (
("00000000000000000000000000000000000000000000000000000000000000000011"),
("00000000000000000000000000000000000000000000000000000111111100001111"),
("00000000000000000000000000000000000000000001111100001111111111001110"),
("00000000000000000000000000001111111100000111111110001111100111001100"),
("00000001110000001111111100001111111110001111001111001100000011001100"),
("11111111100000001111111110011100000111011100000011101100000011001110"),
("11111111100000001100001111011100000111011000000011101100000011001110"),
("00000111000000001100000111011100000111011000000011101100000111000111"),
("00000110000000001100000011011100000111011000000011101111111110000011"),
("00001111000000001100000011011100111110011000000011001111111100000011"),
("00011111110000001100000011011111111100011100000111001100000000000111"),
("00000001110000011100000111011111111000011110011110001100000000011111"),
("00000000110000011100001110011111110000001111111110001100000000011110"),
("00000000111000011111111100011001111000000111111000001100000000000000"),
("00000000110110011111111000011000111100000000000000000000000000000000"),
("00000000110110011111100000000000011110000000000000000000000000000000"),
("01000001110000000000000000000000001110000000000000000000000000000000"),
("11111111100000000000000000000000000100000000000000000000000000000000"),
("11111111000000000000000000000000000000000000000000000000000000000000")
);

----- pitch image
constant pitch_X_size : integer :=68;
constant pitch_Y_size : integer :=15;

--object start
signal X4_begin : integer := 490;
signal Y4_begin : integer := 400;

signal bCoord_X4 : integer := 0;
signal bCoord_Y4 : integer := 0;

signal drawing_X4 : std_logic := '0';
signal drawing_Y4 : std_logic := '0';

type pitch_object is array (0 to pitch_Y_size - 1 , 0 to pitch_X_size - 1) of std_logic;
 constant pitch : pitch_object := (
("00000000000000000000000000000000000000000000000000111110011000000011"),
("00000000000000000000000000000000000111111111100011111110011000000111"),
("00000100001100000000011111100001101111111111100111110000011000000111"),
("00000111001100000001111111110001101111111000000110000000011000000111"),
("00001110011100000001111111111001100000111000001100000000011111111111"),
("00001110011100000011100000011001100000111000001100000000011111111111"),
("00011100011100000011100000011001100000111000011100000000011111110110"),
("00011100011100000011100000011001100000111000011100000000011000000110"),
("00111000011100000011100000111011100000110000001100000000011000000110"),
("00111000011100000011111111110011100000111000001110000000111000000110"),
("01111111111100000011111111100011100000111000001111111100111000000110"),
("01111111111100000011111000000011100000110000000111111100111000000110"),
("11111111111100000011000000000011100000110000000001111000000000000000"),
("00000000011101110011000000000011100000110000000000000000000000000000"),
("00000000011101110011000000000000000000000000000000000000000000000000")
);

begin 

--calculating  x & y coordination for drawing the pictures

-----	

	drawing_X	<= '1' when  (oCoord_X  >=X_begin) and  (oCoord_X < X_begin+flute_X_size) else '0';
	drawing_Y	<= '1' when  (oCoord_Y  >= Y_begin)  and (oCoord_Y  < Y_begin+flute_Y_size) else '0';
            
	bCoord_X   <=  (oCoord_X-X_begin) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y   <= (oCoord_Y-Y_begin) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	
----

	drawing_X2	<= '1' when  (oCoord_X  >=X2_begin) and  (oCoord_X < X2_begin+piano_X_size) else '0';
	drawing_Y2	<= '1' when  (oCoord_Y  >= Y2_begin)  and (oCoord_Y  < Y2_begin+piano_Y_size) else '0';
            
	bCoord_X2   <=  (oCoord_X-X2_begin) when ( drawing_X2 = '1' and  drawing_Y2 = '1'  ) else 0 ; 
	bCoord_Y2   <= (oCoord_Y-Y2_begin) when ( drawing_X2 = '1' and  drawing_Y2 = '1'  ) else 0 ; 
	
-----

	drawing_X3	<= '1' when  (oCoord_X  >=X3_begin) and  (oCoord_X < X3_begin+drop_X_size) else '0';
	drawing_Y3	<= '1' when  (oCoord_Y  >= Y3_begin)  and (oCoord_Y  < Y3_begin+drop_Y_size) else '0';
            
	bCoord_X3   <=  (oCoord_X-X3_begin) when ( drawing_X3 = '1' and  drawing_Y3 = '1'  ) else 0 ; 
	bCoord_Y3   <= (oCoord_Y-Y3_begin) when ( drawing_X3 = '1' and  drawing_Y3 = '1'  ) else 0 ; 
	
-----	
	drawing_X4	<= '1' when  (oCoord_X  >=X4_begin) and  (oCoord_X < X4_begin+pitch_X_size) else '0';
	drawing_Y4	<= '1' when  (oCoord_Y  >= Y4_begin)  and (oCoord_Y  < Y4_begin+pitch_Y_size) else '0';
            
	bCoord_X4   <=  (oCoord_X-X4_begin) when ( drawing_X4 = '1' and  drawing_Y4 = '1'  ) else 0 ; 
	bCoord_Y4   <= (oCoord_Y-Y4_begin) when ( drawing_X4 = '1' and  drawing_Y4 = '1'  ) else 0 ; 
	
process ( RESETn, CLK) 		
 begin 		
	if RESETn = '0' then	
		Pick_inst_request <= '0';
	elsif CLK'event and CLK='1' then
		if  drawing_X='1' and drawing_Y='1' then 
			Pick_inst_request <= flute(bCoord_Y , bCoord_X)  ;
			if  flute_effect = '1' then
				mVGA_RGB <= x"e0" ;-- draw the picture in "red" if it's selected.
			else 
				mVGA_RGB <= x"34" ;-- other wise draw it in "green".
			end if;
		elsif drawing_X2='1' and drawing_Y2='1' then
			Pick_inst_request <= piano(bCoord_Y2 , bCoord_X2);
			if piano_effect = '1' then
				mVGA_RGB <= x"e0" ;
			else 
				mVGA_RGB <= x"34"  ;
			end if;
		elsif drawing_X3='1' and drawing_Y3='1' then
			Pick_inst_request <= drop(bCoord_Y3 , bCoord_X3);
			if drop_effect = '1' then 
				mVGA_RGB <= x"e0" ;
			else 
				mVGA_RGB <= x"34"  ;
			end if;
		elsif drawing_X4='1' and drawing_Y4='1' then
			Pick_inst_request <= pitch(bCoord_Y4 , bCoord_X4);
			if pitch_effect = '1' then
				mVGA_RGB <= x"e0" ;
			else 
				mVGA_RGB <= x"34"  ;
			end if;
		else
			Pick_inst_request <=Notes_screen_request;-- draw the notes on this screen also
			mVGA_RGB <= x"00";
		end if ;
	end if;
end process;
end behav;
library IEEE;
use IEEE.STD_LOGIC_1164.all;

--- drwaing the first screeen
entity Pick_Mode_Screen is
port 	(
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		mVGA_RGB    : out std_logic_vector(7 downto 0);
		Pick_Mode_request	: out std_logic
	);
end Pick_Mode_Screen;

architecture behav of Pick_Mode_Screen is 
--pick size
constant pick_X_size : integer :=90;
constant pick_Y_size : integer :=16;

--object start
signal X_begin : integer := 20;
signal Y_begin : integer := 420 ;

signal bCoord_X : integer := 0;
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';


type pick_object is array (0 to pick_Y_size - 1 , 0 to pick_X_size - 1) of std_logic;
 constant pick: pick_object := (
("000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000"),
("000000000000000000000000000000000000000000000000000000000000010000011111111000111111111000"),
("000000000000000000000000000000000000000000000110000110000011111100011111111100111111100011"),
("000000000000000000000000011000001000000000001110001110000111111110011100011110110000000011"),
("000000000001110001111110011000011100000000001111001111001110000111011000001110110000000000"),
("111111111001110011111110011000111100000000001111011111011100000011011000000110111111100000"),
("111111111101100111000000011001111000000000001111111111011000000011011000000110111111100000"),
("110000011101100110000000111011110000000000011111111011011000000011011000000110110000000000"),
("110000001101101110000000111111100000000000011001110011011000000011011000001110110000000000"),
("110000011101101100000000111111000000000000011001110011011100000111011000011100111011110011"),
("110000111001101110000000111111000000000000011000100011001110011110011111111000111111110011"),
("111111111001101110000000111111100000000000111000100011001111111100011111110000111111110000"),
("111111100001100111000000111001110000000000110000000011000011110000010000000000000000000000"),
("110000000001100111111100110000111000000000110000000011100000000000000000000000000000000000"),
("110000000001100001111100110000011100000000000000000011100000000000000000000000000000000000"),
("110000000001000000000000000000001110000000000000000011100000000000000000000000000000000000")
 );
 


 ----- freeStyle option image
constant freeStyle_X_size : integer :=100;
constant freeStyle_Y_size : integer :=15;

--object start
signal X2_begin : integer := 250;
signal Y2_begin : integer := 400;
 
signal bCoord_X2 : integer := 0;
signal bCoord_Y2 : integer := 0;

signal drawing_X2 : std_logic := '0';
signal drawing_Y2 : std_logic := '0';


type freeStyle_object is array (0 to freeStyle_Y_size - 1 , 0 to freeStyle_X_size - 1) of std_logic;
 constant freeStyle : freeStyle_object := (
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("0011100000000000000001111111000000000000000000000000000000000011111000011000000000000001000000000000"),
("0111100000000000000001111111000000000000000000000000000000000111111000010000000000000001000000000000"),
("0000100000000000000001100000000000000000000000000000000000001100000000111000000000000001000000000000"),
("0000100000000000000001100000011011000111111000011111100000001100000000111110110000011001100011111100"),
("0000100000000000000001111110011100001110011100110001100000000111000000011000011000010001000111001100"),
("0000100000000000000001111110011000001000001101100000110000000011111000011000011000110001000100000110"),
("0000100000000000000001100000011000011111111101111111110000000000011100011000001000100001001111111110"),
("0000100000000000000001100000011000011111111101111111110000000000001100011000001101100001001111111110"),
("0000100000000000000001100000011000001000000001100000000000000000001100011000000111000001000100000000"),
("0001100000000000000001100000011000001110000100110000010000001100011100011000000111000001000111000010"),
("0111111100010000000001100000011000000111111100011111110000001111111000011110000011000001000011111110"),
("0001000000010000000000000000000000000000000000000010000000000000000000000010000010000001000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000")
);


----- Create Tune option image
constant Tune_X_size : integer :=100;
constant Tune_Y_size : integer :=25;

--object start
signal X3_begin : integer := 250;
signal Y3_begin : integer := 430;

signal bCoord_X3 : integer := 0;
signal bCoord_Y3 : integer := 0;

signal drawing_X3 : std_logic := '0';
signal drawing_Y3 : std_logic := '0';

type Tune_object is array (0 to Tune_Y_size - 1 , 0 to Tune_X_size - 1) of std_logic;
 constant Tune : Tune_object := (
("0111110000000000000001111110000000000000000000000000100000000000000001100001100000000000000000000000"),
("0100111000000000000011000010000000000000000000000000100000000000000000100001000000000000000000000000"),
("0000011000000000000110000000011011000111000011110001111000111100000000010011000111100011000100010110"),
("0000011000000000000100000000011110011111110011111001111001111110000000011110001111110011000100011100"),
("0000010000000000000100000000011000010000010000001000100011000011000000001100011000010011000100011000"),
("0000110000000000000100000000011000011111110011111000100011111111000000001100010000011011000100010000"),
("0001100000000000000100000000011000011111110111111000100011111110000000001100011000011011000100010000"),
("0111000000000000000110000000011000011000000110011000100001000000000000001100011000110011001100010000"),
("0111111000100000000011111110011000001111110111111000111001111111000000001100001111110001111100010000"),
("0111111000100000000000011000000000000011000001001000001000001000000000000000000011000000100100010000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000001111100000000000000000000000000001111111110000000000000000000000000000"),
("0000000000000000000000000000011000110000000000000000000000000000000100000000000000000000000000000000"),
("0000000000000000000000000000110000011001100110001000101110000000000100001000110011111000001111000000"),
("0000000000000000000000000000100000011000100110011000110110000000000100001000110011101100111011100000"),
("0000000000000000000000000000100000011000100111011000100011000000000100001000110011000100110000100000"),
("0000000000000000000000000000100000011000101101010000100011000000000100001000110011000100111111100000"),
("0000000000000000000000000000110000011000111001010000100011000000000100001000110011000100110000000000"),
("0000000000000000000000000000111000110000011001110000100011000000000100001000110010000100110000000000"),
("0000000000000000000000000000001111100000011000110000100011000000000100001111110011000100011111100000")
);

----- pro option image
constant pro_X_size : integer :=79;
constant pro_Y_size : integer :=19;

--object start
signal X4_begin : integer := 400;
signal Y4_begin : integer := 415;

signal bCoord_X4 : integer := 0;
signal bCoord_Y4 : integer := 0;

signal drawing_X4 : std_logic := '0';
signal drawing_Y4 : std_logic := '0';

type pro_object is array (0 to pro_Y_size - 1 , 0 to pro_X_size - 1) of std_logic;
 constant pro : pro_object := (
("0000000000000000000000000000000000000000000000000000000000000000000000000000001"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000011"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000011"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000011"),
("0000000000000000000000000000000000000000000000000000001000011111100001111110011"),
("0000000000000000000000000000000000000001100000000011111110011111110011000111011"),
("0111111100000011111100011111100000000011100000000011000110010000010010000011011"),
("0111111100000011111110011000000000000011100000000010000010010000010110000001011"),
("0000011000000010000110010000000000000110110000000010000010010000110110000011011"),
("0000111000000110000110011111000000000110110000000011011110011111100110000011000"),
("0001111100000111111100111111000000001100110000000111111100111111000111000110011"),
("0000001110000111111110110000000000001111111000000110000000110111000011111100011"),
("0000000110000110000110110000000000011111111000000110000000110011100000110000000"),
("0000000110000110011110111111100000011000011000000110000000000001110000000000000"),
("0000000110110111111100111111100000000000001100000000000000000000110000000000000"),
("0100001110100000000000000000000000000000001100000000000000000000000000000000000"),
("1111111100000000000000000000000000000000000000000000000000000000000000000000000"),
("0111111000000000000000000000000000000000000000000000000000000000000000000000000"),
("0001100000000000000000000000000000000000000000000000000000000000000000000000000")
);
begin 


--calculating  x & y coordination for drawing the pictures
-----	

	drawing_X	<= '1' when  (oCoord_X  >=X_begin) and  (oCoord_X < X_begin+pick_X_size) else '0';
	drawing_Y	<= '1' when  (oCoord_Y  >= Y_begin)  and (oCoord_Y  < Y_begin+pick_Y_size) else '0';
            
	bCoord_X   <=  (oCoord_X-X_begin) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y   <= (oCoord_Y-Y_begin) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	
----

	drawing_X2	<= '1' when  (oCoord_X  >=X2_begin) and  (oCoord_X < X2_begin+freeStyle_X_size) else '0';
	drawing_Y2	<= '1' when  (oCoord_Y  >= Y2_begin)  and (oCoord_Y  < Y2_begin+freeStyle_Y_size) else '0';
            
	bCoord_X2   <=  (oCoord_X-X2_begin) when ( drawing_X2 = '1' and  drawing_Y2 = '1'  ) else 0 ; 
	bCoord_Y2   <= (oCoord_Y-Y2_begin) when ( drawing_X2 = '1' and  drawing_Y2 = '1'  ) else 0 ; 
	
-----

	drawing_X3	<= '1' when  (oCoord_X  >=X3_begin) and  (oCoord_X < X3_begin+Tune_X_size) else '0';
	drawing_Y3	<= '1' when  (oCoord_Y  >= Y3_begin)  and (oCoord_Y  < Y3_begin+Tune_Y_size) else '0';
            
	bCoord_X3   <=  (oCoord_X - X3_begin) when ( drawing_X3 = '1' and  drawing_Y3 = '1'  ) else 0 ; 
	bCoord_Y3   <= (oCoord_Y - Y3_begin) when ( drawing_X3 = '1' and  drawing_Y3 = '1'  ) else 0 ; 
	
-----

	drawing_X4	<= '1' when  (oCoord_X  >=X4_begin) and  (oCoord_X < X4_begin+pro_X_size) else '0';
	drawing_Y4	<= '1' when  (oCoord_Y  >= Y4_begin)  and (oCoord_Y  < Y4_begin+pro_Y_size) else '0';
            
	bCoord_X4   <=  (oCoord_X - X4_begin) when ( drawing_X4 = '1' and  drawing_Y4 = '1'  ) else 0 ; 
	bCoord_Y4   <= (oCoord_Y - Y4_begin) when ( drawing_X4 = '1' and  drawing_Y4 = '1'  ) else 0 ; 	
process ( RESETn, CLK) 		
 begin
   	mVGA_RGB <= x"6F" ;	
	if RESETn = '0' then	
		Pick_Mode_request <= '0';
	elsif CLK'event and CLK='1' then
		if  drawing_X = '1'  and drawing_Y = '1'  then 
			Pick_Mode_request <= pick(bCoord_Y , bCoord_X)  ;
		elsif drawing_X2 = '1'  and drawing_Y2 = '1'  then
			Pick_Mode_request <= freeStyle(bCoord_Y2 , bCoord_X2);
		elsif drawing_X4 = '1'  and drawing_Y4 = '1'  then
			Pick_Mode_request <= pro(bCoord_Y4 , bCoord_X4);
		else 
			Pick_Mode_request <= drawing_X3 and drawing_Y3 and Tune(bCoord_Y3 , bCoord_X3);
		end if ;
	end if;
end process;
end behav;
constant_0_inst : constant_0 PORT MAP (
		result	 => result_sig
	);
